* C:\FOSSEE\eSim\library\SubcircuitLibrary\HA_kalyan\HA_kalyan.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 10/02/22 12:57:29

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
X2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad4_ xor_gate_kalyan		
X1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ and_kalyan		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ PORT		

.end
